
.MODEL MBRB1645 D (IS=500N N=1.18295 BV=51 IBV=10M RS=5.9528M CJO=3.23313N VJ=700M
M=493.226M EG=900M XTI=2 RL=875.289K T_MEASURED=25°C)
